module reg_file(
    input clk,
    input we,                   // write enable
    input [4:0] ra1, ra2, rw,   // read addresses 1, 2 and write address
    input [31:0] wd,            // write data
    output [31:0] rd1, rd2      // read data 1, read data 2
);

    reg [31:0] regs [31:0];

    assign rd1 = (ra1 == 0) ? 32'b0 : regs[ra1];
    assign rd2 = (ra2 == 0) ? 32'b0 : regs[ra2];

    always @(posedge clk) begin
        regs[0] <= 32'b0;   // enforce $zero
        if (we && (rw != 0))
            regs[rw] <= wd;
    end
endmodule
